// Author: Graham Nygard, Robert Wagner

module IFID_reg(clk, )

//INPUTS
input clk;

//OUTPUTS


always @(posedge clk) begin
	q <= d;
end

endmodule