// Author: Graham Nygard, Robert Wagner

module WB_Unit(clk, 
	mem_read_data_in, reg_rd_in, ret_future_in, alu_result_in
	)

//INPUTS
input clk;
input mem_read_data_in;
input reg_rd_in;
input ret_future_in;
input alu_result_in;

//OUTPUTS


//MODULE INSTANTIATIONS



endmodule