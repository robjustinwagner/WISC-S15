
module WISC_S15_top_level ( clk, rst );
  input clk, rst;


endmodule

