// Author: Graham Nygard, Robert Wagner

module Sign_Ext_Unit(arith_imm_in, load_save_imm_in,
                     sign_ext);
