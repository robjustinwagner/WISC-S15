// Author: Graham Nygard, Robert Wagner

module WB_Unit(clk, );

//INPUTS
input clk;

//OUTPUTS


//MODULE INSTANTIATIONS



endmodule