// Author: Graham Nygard, Robert Wagner

module MEMWB_reg(clk, )

//INPUTS
input clk;

//OUTPUTS


always @(posedge clk) begin
	q <= d;
end

endmodule