// Author: Graham Nygard, Robert Wagner

module HDT_Unit();
