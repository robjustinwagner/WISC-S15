// Author: Graham Nygard, Robert Wagner

module EXMEM_reg(clk, )

//INPUTS
input clk;

//OUTPUTS


always @(posedge clk) begin
	q <= d;
end

endmodule